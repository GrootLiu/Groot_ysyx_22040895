`include "../include/include.v"

module sext (input wire rst,
             input wire immsel_i_sext,
             input wire[`imm1Length] imm1_i_sext,
             input wire[`imm2Length] imm1_i_sext,
             output wire[`RegBus] simm_o_sext);

    
    
    
endmodule //sext
